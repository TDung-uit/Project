module shift1R(I,O);
input [4:0] I;
output [4:0] O;
	assign O = I >> 1;

endmodule
